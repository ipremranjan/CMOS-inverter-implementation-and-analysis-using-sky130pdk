magic
tech sky130A
timestamp 1705035004
<< nwell >>
rect -150 -50 150 370
<< nmos >>
rect -10 -200 5 -100
<< pmos >>
rect -10 -5 5 205
<< ndiff >>
rect -50 -110 -10 -100
rect -50 -190 -40 -110
rect -20 -190 -10 -110
rect -50 -200 -10 -190
rect 5 -110 50 -100
rect 5 -190 20 -110
rect 40 -190 50 -110
rect 5 -200 50 -190
<< pdiff >>
rect -60 195 -10 205
rect -60 5 -50 195
rect -25 5 -10 195
rect -60 -5 -10 5
rect 5 195 55 205
rect 5 5 20 195
rect 45 5 55 195
rect 5 -5 55 5
<< ndiffc >>
rect -40 -190 -20 -110
rect 20 -190 40 -110
<< pdiffc >>
rect -50 5 -25 195
rect 20 5 45 195
<< psubdiff >>
rect -65 -240 70 -230
rect -65 -260 -50 -240
rect 50 -260 70 -240
rect -65 -275 70 -260
<< nsubdiff >>
rect -85 315 70 325
rect -85 285 -70 315
rect 55 285 70 315
rect -85 275 70 285
<< psubdiffcont >>
rect -50 -260 50 -240
<< nsubdiffcont >>
rect -70 285 55 315
<< poly >>
rect -10 205 5 260
rect -10 -30 5 -5
rect -60 -40 5 -30
rect -60 -60 -50 -40
rect -25 -60 5 -40
rect -60 -70 5 -60
rect 65 -40 110 -30
rect 65 -60 75 -40
rect 100 -60 110 -40
rect 65 -70 110 -60
rect -10 -100 5 -70
rect -10 -215 5 -200
<< polycont >>
rect -50 -60 -25 -40
rect 75 -60 100 -40
<< locali >>
rect -85 320 70 325
rect -85 315 -40 320
rect 35 315 70 320
rect -85 285 -70 315
rect 55 285 70 315
rect -85 280 -40 285
rect 35 280 70 285
rect -85 275 70 280
rect -60 195 -15 275
rect -60 5 -50 195
rect -25 5 -15 195
rect -60 -5 -15 5
rect 10 195 55 205
rect 10 5 20 195
rect 45 5 55 195
rect 10 -5 55 5
rect 15 -30 50 -5
rect -60 -40 -15 -30
rect -60 -60 -50 -40
rect -25 -60 -15 -40
rect -60 -70 -15 -60
rect 15 -40 110 -30
rect 15 -60 75 -40
rect 100 -60 110 -40
rect 15 -70 110 -60
rect 15 -100 50 -70
rect -50 -110 -15 -100
rect -50 -190 -40 -110
rect -20 -190 -15 -110
rect -50 -230 -15 -190
rect 10 -110 50 -100
rect 10 -190 20 -110
rect 40 -190 50 -110
rect 10 -200 50 -190
rect -65 -235 70 -230
rect -65 -240 -30 -235
rect 30 -240 70 -235
rect -65 -260 -50 -240
rect 50 -260 70 -240
rect -65 -270 -30 -260
rect 30 -270 70 -260
rect -65 -275 70 -270
<< viali >>
rect -40 315 35 320
rect -40 285 35 315
rect -40 280 35 285
rect -50 -60 -25 -40
rect 75 -60 100 -40
rect -30 -240 30 -235
rect -30 -260 30 -240
rect -30 -270 30 -260
<< metal1 >>
rect -280 320 330 325
rect -280 280 -40 320
rect 35 280 330 320
rect -280 275 330 280
rect -270 -40 -15 -30
rect -270 -60 -50 -40
rect -25 -60 -15 -40
rect -270 -70 -15 -60
rect 15 -40 330 -30
rect 15 -60 75 -40
rect 100 -60 330 -40
rect 15 -70 330 -60
rect -270 -235 330 -230
rect -270 -270 -30 -235
rect 30 -270 330 -235
rect -270 -275 330 -270
<< labels >>
rlabel metal1 250 295 250 295 1 vdd
rlabel metal1 230 -250 230 -250 1 vss
rlabel metal1 275 -55 290 -40 1 out
rlabel metal1 -255 -60 -235 -40 1 in
<< end >>
